module sr_latch(
    input s, r,
    output q, qb
);
nand u1 (q, s, qb);
nand u2 (qb, r, q);

endmodule
